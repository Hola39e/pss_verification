package pss_vseq_lib_pkg;

    import uvm_pkg::*;
    `include "uvm_macros.svh"
    
    import ahb_agent_pkg::*;
    import spi_agent_pkg::*;
    import gpio_agent_pkg::*;
    import gpio_bus_sequence_lib_pkg::*;
    import gpio_sequence_lib_pkg::*;
    import spi_bus_sequence_lib_pkg::*;
    import spi_sequence_lib_pkg::*;
    import pss_env_pkg::*;
    
    `include "bridge_basic_rw_vseq.svh"
    `include "pss_vseq_base.svh"
    `include "gpio_outputs_vseq.svh"
    `include "spi_interrupt_vseq.svh"
    `include "spi_polling_vseq.svh"
    
    
    endpackage: pss_vseq_lib_pkg