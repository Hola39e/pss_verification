package gpio_test_lib_pkg;

    // Standard UVM import & include:
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    
    // Any further package imports:
    import gpio_env_pkg::*;
    import apb_agent_pkg::*;
    import gpio_agent_pkg::*;
    import gpio_register_pkg::*;
    import gpio_virtual_sequence_lib_pkg::*;
    import register_layering_pkg::*;
    
    // Includes:
    `include "gpio_test_base.svh"
    `include "gpio_input_test.svh"
    
    endpackage: gpio_test_lib_pkg
    