
package pss_test_lib_pkg;

    // Standard UVM import & include:
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    
    // Any further package imports:
    import spi_env_pkg::*;
    import apb_agent_pkg::*;
    import ahb_agent_pkg::*;
    import spi_agent_pkg::*;
    import gpio_agent_pkg::*;
    import gpio_env_pkg::*;
    import pss_env_pkg::*;
    import pss_vseq_lib_pkg::*;
	import gpio_register_model_pkg::*;
	import spi_reg_pkg::*;
	import pss_register_model_pkg::*;
	
    
    // Includes:
    `include "pss_test_base.svh"
    // `include "pss_test.svh"
    // `include "pss_gpio_outputs_test.svh"
    // `include "pss_spi_polling_test.svh"
    // `include "pss_spi_interrupt_test.svh"
    
    endpackage: pss_test_lib_pkg
    