package apb_agent_pkg;
    import uvm_pkg::*;
	
	import register_layering_pkg::*;
	
    `include "uvm_macros.svh"
    `include "apb_seq_item.svh"
    `include "apb_agent_config.svh"
    `include "apb_driver.svh"
    `include "apb_coverage_monitor.svh"
    `include "apb_monitor.svh"
    `include "apb_sequencer.svh"
    `include "apb_agent.svh"

    // Utility Sequences
    `include "apb_seq.svh"
    `include "apb_read_seq.svh"
    `include "apb_write_seq.svh"
    `include "apb_register_adapter.svh"
    `include "apb2reg_adapter.sv"
endpackage
