interface spi_if;

  logic clk;
  logic[7:0] cs;
  logic miso;
  logic mosi;
endinterface: spi_if
