package gpio_agent_pkg;

    import uvm_pkg::*;

    `include "uvm_marcos.svh"

    `include "gpio_seq_item.svh"
    `include "gpio_agent_config.svh"
    `include "gpio_driver.svh"
    `include "gpio_monitor.svh"
    `include "gpio_sequencer.svh"
    `include "gpio_agent.svh"

    // Utility Sequences
    `include "gpio_seq.svh"
endpackage