interface serial_if;
    logic sdata;
    logic clk;
endinterface