class gpio_output_vseq extends pss_vseq_base;

    `uvm_object_utils(gpio_output_vseq)

    function new(string name = "gpio_outputs_vseq");
        super.new(name);
    endfunction

    task body;
        // -----------------need to change
    endtask

endclass