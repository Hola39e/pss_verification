interface intr_if;
    logic IRQ;
endinterface