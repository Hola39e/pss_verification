
package gpio_rgm_test_lib_pkg;

    // Standard UVM import & include:
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    
    // Any further package imports:
    import gpio_env_pkg::*;
    import apb_agent_pkg::*;
    import gpio_agent_pkg::*;
    import gpio_register_model_pkg::*;
    import gpio_rgm_virtual_sequence_pkg::*;
	
    
    // Includes:
    `include "gpio_rgm_test_base.sv"
    `include "gpio_rgm_input_test.sv"
    `include "gpio_rgm_input_read_test.sv"
endpackage: gpio_rgm_test_lib_pkg
    