package spi_agent_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"

//import spi_register_pkg::*;

`include "spi_seq_item.svh"
`include "spi_agent_config.svh"
`include "spi_driver.svh"
`include "spi_monitor.svh"
`include "spi_sequencer.svh"
`include "spi_agent.svh"

// Utility Sequences
`include "spi_seq.svh"

endpackage: spi_agent_pkg