package pss_env_pkg;

// Standard UVM import & include:
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    import gpio_env_pkg::*;
    import spi_env_pkg::*;
    import ahb_agent_pkg::*;
    import spi_agent_pkg::*;
    import gpio_agent_pkg::*;
    `include "pss_env_config.svh"
    `include "pss_virtual_sequencer.svh"
    `include "pss_env.svh"
    
endpackage: pss_env_pkg
